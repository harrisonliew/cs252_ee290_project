../../../../../../Verilog HD Sensor Fusion/const.vh